module uncodeable
  #(
    P = 0
    )
   (
    input logic clk,
    input logic rst,
    );

endmodule
